class pd_debug_cascade_test extends pd_debug_base_test;
    `uvm_component_utils(pd_debug_cascade_test)

    pd_debug_cascade_sequence cascade_seq;

    function new(string name = "pd_debug_cascade_test", uvm_component parent = null);
            super.new(name, parent);
        endfunction 


    // virtual function void build_phase(uvm_phase phase);
    //     super.build_phase(phase);

    //     pd_debug_agt_cfg.driving_cycles = 2;

    // endfunction

    virtual task run_phase(uvm_phase phase);
        super.run_phase(phase);

        cascade_seq = pd_debug_cascade_sequence::type_id::create("cascade_seq");

        phase.raise_objection(this, get_type_name());

        //main_sequence
        `uvm_info(get_type_name(), "Stimulus Generation Started", UVM_LOW);

        //Match Sequence
        `uvm_info(get_type_name(), "Cascade Sequence Started \n", UVM_LOW);
        cascade_seq.init_start(pd_debug_agt_cfg.pd_debug_sqr);
        `uvm_info(get_type_name(), "Cascade Sequence Ended \n", UVM_LOW);

        `uvm_info(get_type_name(), "Stimulus Generation Ended", UVM_LOW);

        phase.drop_objection(this, get_type_name());
        
    endtask
endclass